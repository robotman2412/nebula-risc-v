`ifndef AHB_LITE_UVC_ENV_TOP_PKG
`define AHB_LITE_UVC_ENV_TOP_PKG

package ahb_lite_uvc_env_top_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

import ahb_lite_uvc_pkg::*;

`include "ahb_lite_uvc_cfg_top.sv"
`include "ahb_lite_uvc_env_top.sv"

endpackage : ahb_lite_uvc_env_top_pkg

`endif // AHB_LITE_UVC_ENV_TOP_PKG
