`ifndef AHB_LITE_UVC_PKG_SV
`define AHB_LITE_UVC_PKG_SV

package ahb_lite_uvc_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ahb_lite_uvc_common.sv"
`include "ahb_lite_uvc_item.sv"
`include "ahb_lite_uvc_seq_lib.sv"
`include "ahb_lite_uvc_agent_cfg.sv"
`include "ahb_lite_uvc_driver.sv"
`include "ahb_lite_uvc_sequencer.sv"
`include "ahb_lite_uvc_monitor.sv"
`include "ahb_lite_uvc_subscriber.sv"
`include "ahb_lite_uvc_agent.sv"
`include "ahb_lite_uvc_env_cfg.sv"
`include "ahb_lite_uvc_env.sv"

endpackage : ahb_lite_uvc_pkg

`include "ahb_lite_uvc_if.sv"

`endif // VENV_UVC_PKG_SV
